emoncore
R7 5 11 22
R13 9 14 100k
R1 6 7 22k
R4 2 11 22
R11 10 1 4.7k
C1 0 7 1µF IC=0
R9 17 11 22
R3 3 11 22
R10 8 1 4.7k
R2 0 7 22k
R8 13 11 22
R14 11 14 10k
R5 4 11 22
R6 16 11 22
R12 15 0 220

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
